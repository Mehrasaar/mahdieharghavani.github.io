** Profile: "SCHEMATIC1-Example 2 Simulation"  [ C:\USERS\ASUS\PSpice Projects\example 2 simulation-SCHEMATIC1-Example 2 Simulation.sim ] 

** Creating circuit file "example 2 simulation-SCHEMATIC1-Example 2 Simulation.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\example 2 simulation-SCHEMATIC1.net" 


.END
