** Profile: "SCHEMATIC1-Simulation1"  [ C:\USERS\ASUS\PSpice Projects\bias point simulations-SCHEMATIC1-Simulation1.sim ] 

** Creating circuit file "bias point simulations-SCHEMATIC1-Simulation1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 0.01 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\bias point simulations-SCHEMATIC1.net" 


.END
